module carry_flag (input sel, cout, output flag);

and n1(flag,sel,cout);

endmodule 