module OR_Gate(input a,b,
				output s);	
or n1(s,a,b);
endmodule
