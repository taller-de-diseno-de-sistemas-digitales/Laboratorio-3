module XOR_Gate(input a,b,
				output s);	
xor n1(s,a,b);
endmodule

