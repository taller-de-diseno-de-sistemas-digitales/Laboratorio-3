module NOT_Gate(input a,
				output s);	
not n1(s,a);
endmodule
