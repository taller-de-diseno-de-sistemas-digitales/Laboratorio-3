module AND_Gate(input a,b,
				output s);	
and n1(s,a,b);
endmodule
