module negative_flag (input in, output flag);

not n1(flag,~in);

endmodule 